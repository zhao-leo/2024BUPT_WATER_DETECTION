`timescale 1ns/1ps
module water_detection_test;
reg clk;
reg btn7;
reg btn0;
reg [3:0] row_in;
wire [7:0] row;
wire [6:0] segment7;
wire [3:0] col;
wire [7:0] green_led;
wire [7:0] red_led;
wire [7:0] select ;
wire beep;
wire dp;
water_detection water_detection1(
    .clk(clk),
    .btn7(btn7),
    .btn0(btn0),
    .row_in(row_in),
    .segment7(segment7),
    .select(select),
    .col(col),
    .row(row),
    .green_led(green_led),
    .red_led(red_led),
    .beep(beep),
    .dp(dp)
);
initial begin
    clk = 1'b0;
    btn7 = 1'b0;
    btn0 = 1'b0;
    row_in = 4'b1111;
    forever #50 clk = ~clk;
end
initial begin
    #100;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;

    #1500;

    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;
    row_in = 4'b1011;
    #100;
    row_in = 4'b1111;
    #300;

    #1500;
    btn0 = 1'b1;
    #2000;
    btn0 = 1'b0;
    #1000;
    btn7 = 1'b1;
    #2000;
    btn7 = 1'b0;
    #1000;
    #10000;
    btn0 = 1'b1;
    #2000;
    btn0 = 1'b0;
    #1000;


    $finish;

end

initial begin
    $dumpfile("tb_water_detection.vcd");
    $dumpvars(0,water_detection_test);
end
endmodule